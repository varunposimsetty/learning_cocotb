module ifc_or(
    input CLK
);
endmodule